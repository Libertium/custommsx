-- 
-- SlotCounter.vhd 
--
-- Copyright (c) 2006 Mitsutaka Okazaki (brezza@pokipoki.org)
-- All rights reserved.
-- 
-- Redistribution and use of this source code or any derivative works, are 
-- permitted provided that the following conditions are met:
--
-- 1. Redistributions of source code must retain the above copyright notice, 
--    this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright 
--    notice, this list of conditions and the following disclaimer in the 
--    documentation and/or other materials provided with the distribution.
-- 3. Redistributions may not be sold, nor may they be used in a commercial 
--    product or activity without specific prior written permission.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS 
-- "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED 
-- TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR 
-- PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR 
-- CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, 
-- EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, 
-- PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
-- OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, 
-- WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR 
-- OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF 
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--
--

--
--	modified by t.hara
--

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;

entity SlotCounter is 
	generic (
		delay	: integer
	);
	port (
		clk		: in	std_logic;
		reset	: in	std_logic;
		clkena	: in	std_logic;

		slot	: out	std_logic_vector( 4 downto 0 );
		stage	: out	std_logic_vector( 1 downto 0 )
	);
end SlotCounter;

architecture rtl of SlotCounter is
	signal ff_count		: std_logic_vector( 6 downto 0 );
begin

	process( reset, clk )
	begin
		if( reset = '1' )then
			ff_count <= "1000111" - delay;
		elsif( clk'event and clk='1' )then
			if( clkena ='1' )then
				if( ff_count = "1000111" )then		-- 71
					ff_count <= (others => '0');
				else
					ff_count <= ff_count + 1;
				end if;
			end if;
		end if;
	end process;

	stage	<= ff_count( 1 downto 0 );		--	0�`3 �ŏz�� 
	slot	<= ff_count( 6 downto 2 );		--	0�`17 �ŏz�� 
end rtl;
